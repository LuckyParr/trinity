module backend (
    input wire               clock,
    input wire               rst_n,
    input wire [`LREG_RANGE] rs1,
    input wire [`LREG_RANGE] rs2,
    input wire [`LREG_RANGE] rd,
    input wire [ `SRC_RANGE] src1,
    input wire [ `SRC_RANGE] src2,
    input wire [ `SRC_RANGE] imm,
    input wire               src1_is_reg,
    input wire               src2_is_reg,
    input wire               need_to_wb,

    //sig below is control transfer(xfer) type
    input wire [    `CX_TYPE_RANGE] cx_type,
    input wire                      is_unsigned,
    input wire [   `ALU_TYPE_RANGE] alu_type,
    input wire                      is_word,
    input wire                      is_load,
    input wire                      is_imm,
    input wire                      is_store,
    input wire [               3:0] ls_size,
    input wire [`MULDIV_TYPE_RANGE] muldiv_type,
    input wire [         `PC_RANGE] pc,
    input wire [      `INSTR_RANGE] instr,

    //write back lreg 
    output wire                 wb_valid,
    output wire [`RESULT_RANGE] wb_data

);
    exu u_exu (
        .rs1            (rs1),
        .rs2            (rs2),
        .rd             (rd),
        .src1           (src1),
        .src2           (src2),
        .imm            (imm),
        .src1_is_reg    (src1_is_reg),
        .src2_is_reg    (src2_is_reg),
        .need_to_wb     (need_to_wb),
        .cx_type        (cx_type),
        .is_unsigned    (is_unsigned),
        .alu_type       (alu_type),
        .is_word        (is_word),
        .is_load        (is_load),
        .is_imm         (is_imm),
        .is_store       (is_store),
        .ls_size        (ls_size),
        .muldiv_type    (muldiv_type),
        .pc             (pc),
        .instr          (instr),
        .redirect_valid (redirect_valid),
        .redirect_target(redirect_target),
        .ls_address     (ls_address),
        .alu_result     (alu_result),
        .bju_result     (bju_result),
        .muldiv_result  (muldiv_result)
    );

    exu_mem_reg u_exu_mem_reg (
        .clock            (clock),
        .rst_n            (rst_n),
        .stall             ()
        .rs1              (rs1),
        .rs2              (rs2),
        .rd               (rd),
        .src1             (src1),
        .src2             (src2),
        .imm              (imm),
        .src1_is_reg      (src1_is_reg),
        .src2_is_reg      (src2_is_reg),
        .need_to_wb       (need_to_wb),
        .cx_type          (cx_type),
        .is_unsigned      (is_unsigned),
        .alu_type         (alu_type),
        .is_word          (is_word),
        .is_load          (is_load),
        .is_imm           (is_imm),
        .is_store         (is_store),
        .ls_size          (ls_size),
        .muldiv_type      (muldiv_type),
        .pc               (pc),
        .instr            (instr),
        .ls_address       (ls_address),
        .alu_result       (alu_result),
        .bju_result       (bju_result),
        .muldiv_result    (muldiv_result),
        .out_rs1          (mem_rs1),
        .out_rs2          (mem_rs2),
        .out_rd           (mem_rd),
        .out_src1         (mem_src1),
        .out_src2         (mem_src2),
        .out_imm          (mem_imm),
        .out_src1_is_reg  (mem_src1_is_reg),
        .out_src2_is_reg  (mem_src2_is_reg),
        .out_need_to_wb   (mem_need_to_wb),
        .out_cx_type      (mem_cx_type),
        .out_is_unsigned  (mem_is_unsigned),
        .out_alu_type     (mem_alu_type),
        .out_is_word      (mem_is_word),
        .out_is_load      (mem_is_load),
        .out_is_imm       (mem_is_imm),
        .out_is_store     (mem_is_store),
        .out_ls_size      (mem_ls_size),
        .out_muldiv_type  (mem_muldiv_type),
        .out_pc           (mem_pc),
        .out_instr        (mem_instr),
        .out_ls_address   (mem_ls_address),
        .out_alu_result   (mem_alu_result),
        .out_bju_result   (mem_bju_result),
        .out_muldiv_result(mem_muldiv_result)
    );

    mem u_mem (
        .clock        (clock),
        .rst_n        (rst_n),
        .is_load      (mem_is_load),
        .is_store     (mem_is_store),
        .src2         (mem_src2),
        .ls_address   (mem_ls_address),
        .ls_size      (mem_ls_size),
        .read_valid   (read_valid),
        .read_ready   (read_ready),
        .read_address (read_address),
        .read_done    (read_done),
        .read_data    (read_data),
        .write_valid  (write_valid),
        .write_ready  (write_ready),
        .write_address(write_address),
        .write_data   (write_data),
        .write_mask   (write_mask),
        .write_done   (write_done)
    );


    exu_mem_reg u_mem_wb_reg (
        .clock            (clock),
        .rst_n            (rst_n),
        .stall          (1'b0),
        .rs1              (mem_rs1),
        .rs2              (mem_rs2),
        .rd               (mem_rd),
        .src1             (mem_src1),
        .src2             (mem_src2),
        .imm              (mem_imm),
        .src1_is_reg      (mem_src1_is_reg),
        .src2_is_reg      (mem_src2_is_reg),
        .need_to_wb       (mem_need_to_wb),
        .cx_type          (mem_cx_type),
        .is_unsigned      (mem_is_unsigned),
        .alu_type         (mem_alu_type),
        .is_word          (mem_is_word),
        .is_load          (mem_is_load),
        .is_imm           (mem_is_imm),
        .is_store         (mem_is_store),
        .ls_size          (mem_ls_size),
        .muldiv_type      (mem_muldiv_type),
        .pc               (mem_pc),
        .instr            (mem_instr),
        .ls_address       (mem_ls_address),
        .alu_result       (mem_alu_result),
        .bju_result       (mem_bju_result),
        .muldiv_result    (mem_muldiv_result),
        .out_rs1          (out_rs1),
        .out_rs2          (out_rs2),
        .out_rd           (out_rd),
        .out_src1         (out_src1),
        .out_src2         (out_src2),
        .out_imm          (out_imm),
        .out_src1_is_reg  (out_src1_is_reg),
        .out_src2_is_reg  (out_src2_is_reg),
        .out_need_to_wb   (out_need_to_wb),
        .out_cx_type      (out_cx_type),
        .out_is_unsigned  (out_is_unsigned),
        .out_alu_type     (out_alu_type),
        .out_is_word      (out_is_word),
        .out_is_load      (out_is_load),
        .out_is_imm       (out_is_imm),
        .out_is_store     (out_is_store),
        .out_ls_size      (out_ls_size),
        .out_muldiv_type  (out_muldiv_type),
        .out_pc           (out_pc),
        .out_instr        (out_instr),
        .out_ls_address   (out_ls_address),
        .out_alu_result   (out_alu_result),
        .out_bju_result   (out_bju_result),
        .out_muldiv_result(out_muldiv_result)
    );



    wire commit_valid = out_alu_type | out_cx_type | out_muldiv_type | is_load | is_store;
    DifftestInstrCommit u_DifftestInstrCommit (
        .clock     (clock),
        .enable    (1'b1),
        .io_valid  (commit_valid),
        .io_skip   (1'b0),
        .io_isRVC  (1'b0),
        .io_rfwen  (out_need_to_wb),
        .io_fpwen  (1'b0),
        .io_vecwen (1'b0),
        .io_wpdest (out_rd),
        .io_wdest  (out_rd),
        .io_pc     (out_pc),
        .io_instr  (out_instr),
        .io_robIdx ('b0),
        .io_lqIdx  ('b0),
        .io_sqIdx  ('b0),
        .io_isLoad ('b0),
        .io_isStore('b0),
        .io_nFused ('b0),
        .io_special('b0),
        .io_coreid ('b0),
        .io_index  ('b0)
    );
endmodule
