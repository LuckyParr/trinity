
module DifftestArchVecRegState(
  input         clock,
  input         enable,
  input  [63:0] io_value_0,
  input  [63:0] io_value_1,
  input  [63:0] io_value_2,
  input  [63:0] io_value_3,
  input  [63:0] io_value_4,
  input  [63:0] io_value_5,
  input  [63:0] io_value_6,
  input  [63:0] io_value_7,
  input  [63:0] io_value_8,
  input  [63:0] io_value_9,
  input  [63:0] io_value_10,
  input  [63:0] io_value_11,
  input  [63:0] io_value_12,
  input  [63:0] io_value_13,
  input  [63:0] io_value_14,
  input  [63:0] io_value_15,
  input  [63:0] io_value_16,
  input  [63:0] io_value_17,
  input  [63:0] io_value_18,
  input  [63:0] io_value_19,
  input  [63:0] io_value_20,
  input  [63:0] io_value_21,
  input  [63:0] io_value_22,
  input  [63:0] io_value_23,
  input  [63:0] io_value_24,
  input  [63:0] io_value_25,
  input  [63:0] io_value_26,
  input  [63:0] io_value_27,
  input  [63:0] io_value_28,
  input  [63:0] io_value_29,
  input  [63:0] io_value_30,
  input  [63:0] io_value_31,
  input  [63:0] io_value_32,
  input  [63:0] io_value_33,
  input  [63:0] io_value_34,
  input  [63:0] io_value_35,
  input  [63:0] io_value_36,
  input  [63:0] io_value_37,
  input  [63:0] io_value_38,
  input  [63:0] io_value_39,
  input  [63:0] io_value_40,
  input  [63:0] io_value_41,
  input  [63:0] io_value_42,
  input  [63:0] io_value_43,
  input  [63:0] io_value_44,
  input  [63:0] io_value_45,
  input  [63:0] io_value_46,
  input  [63:0] io_value_47,
  input  [63:0] io_value_48,
  input  [63:0] io_value_49,
  input  [63:0] io_value_50,
  input  [63:0] io_value_51,
  input  [63:0] io_value_52,
  input  [63:0] io_value_53,
  input  [63:0] io_value_54,
  input  [63:0] io_value_55,
  input  [63:0] io_value_56,
  input  [63:0] io_value_57,
  input  [63:0] io_value_58,
  input  [63:0] io_value_59,
  input  [63:0] io_value_60,
  input  [63:0] io_value_61,
  input  [63:0] io_value_62,
  input  [63:0] io_value_63,
  input  [ 7:0] io_coreid
);
`ifndef SYNTHESIS
`ifdef DIFFTEST

import "DPI-C" function void v_difftest_ArchVecRegState (
  input   longint io_value_0,
  input   longint io_value_1,
  input   longint io_value_2,
  input   longint io_value_3,
  input   longint io_value_4,
  input   longint io_value_5,
  input   longint io_value_6,
  input   longint io_value_7,
  input   longint io_value_8,
  input   longint io_value_9,
  input   longint io_value_10,
  input   longint io_value_11,
  input   longint io_value_12,
  input   longint io_value_13,
  input   longint io_value_14,
  input   longint io_value_15,
  input   longint io_value_16,
  input   longint io_value_17,
  input   longint io_value_18,
  input   longint io_value_19,
  input   longint io_value_20,
  input   longint io_value_21,
  input   longint io_value_22,
  input   longint io_value_23,
  input   longint io_value_24,
  input   longint io_value_25,
  input   longint io_value_26,
  input   longint io_value_27,
  input   longint io_value_28,
  input   longint io_value_29,
  input   longint io_value_30,
  input   longint io_value_31,
  input   longint io_value_32,
  input   longint io_value_33,
  input   longint io_value_34,
  input   longint io_value_35,
  input   longint io_value_36,
  input   longint io_value_37,
  input   longint io_value_38,
  input   longint io_value_39,
  input   longint io_value_40,
  input   longint io_value_41,
  input   longint io_value_42,
  input   longint io_value_43,
  input   longint io_value_44,
  input   longint io_value_45,
  input   longint io_value_46,
  input   longint io_value_47,
  input   longint io_value_48,
  input   longint io_value_49,
  input   longint io_value_50,
  input   longint io_value_51,
  input   longint io_value_52,
  input   longint io_value_53,
  input   longint io_value_54,
  input   longint io_value_55,
  input   longint io_value_56,
  input   longint io_value_57,
  input   longint io_value_58,
  input   longint io_value_59,
  input   longint io_value_60,
  input   longint io_value_61,
  input   longint io_value_62,
  input   longint io_value_63,
  input      byte io_coreid
);


  always @(posedge clock) begin
    if (enable)
      v_difftest_ArchVecRegState (io_value_0, io_value_1, io_value_2, io_value_3, io_value_4, io_value_5, io_value_6, io_value_7, io_value_8, io_value_9, io_value_10, io_value_11, io_value_12, io_value_13, io_value_14, io_value_15, io_value_16, io_value_17, io_value_18, io_value_19, io_value_20, io_value_21, io_value_22, io_value_23, io_value_24, io_value_25, io_value_26, io_value_27, io_value_28, io_value_29, io_value_30, io_value_31, io_value_32, io_value_33, io_value_34, io_value_35, io_value_36, io_value_37, io_value_38, io_value_39, io_value_40, io_value_41, io_value_42, io_value_43, io_value_44, io_value_45, io_value_46, io_value_47, io_value_48, io_value_49, io_value_50, io_value_51, io_value_52, io_value_53, io_value_54, io_value_55, io_value_56, io_value_57, io_value_58, io_value_59, io_value_60, io_value_61, io_value_62, io_value_63, io_coreid);
  end
`endif
`endif
endmodule
