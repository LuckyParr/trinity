module #()
(

);

/* --------------------- write instr0 and instr1 to rob --------------------- */


/* ------- read instr0 and instr1 rs1 rs2 busy status from busy_vector ------ */

/* ------- check if instr1 need to sleep due to raw hazard with instr0 ------ */

/* ------------------------------ set sleep bit ----------------------------- */

/* ------------- send instr0 instr1 and sleep bit to issue queue ------------ */




endmodule