// `include "deinfes.sv"
// module writeback (
//     input wire [`LREG_RANGE] rd,
//     input wire [`RESULT_RANGE] write_back_value,
//     input wire need_to_wb,


// );
    
// endmodule