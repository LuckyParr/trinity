module #()
(

);
//issue queue is a 2d reg array
/* ------------------- use findfirst_2availableblock to get place to enqueue 2 instr at same time ------------------- */



/* ---------- receive writeback info to wakeup instr in issue queue --------- */



/* ---------------- use findfirst to find first non-sleep instr to send to fu --------------- */




/* ------------------ get reg content from physical regfile ----------------- */




/* ---------------------------- send instr to fu ---------------------------- */





endmodule