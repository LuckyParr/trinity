
module DifftestSbufferEvent(
  input         clock,
  input         enable,
  input         io_valid,
  input  [63:0] io_addr,
  input  [ 7:0] io_data_0,
  input  [ 7:0] io_data_1,
  input  [ 7:0] io_data_2,
  input  [ 7:0] io_data_3,
  input  [ 7:0] io_data_4,
  input  [ 7:0] io_data_5,
  input  [ 7:0] io_data_6,
  input  [ 7:0] io_data_7,
  input  [ 7:0] io_data_8,
  input  [ 7:0] io_data_9,
  input  [ 7:0] io_data_10,
  input  [ 7:0] io_data_11,
  input  [ 7:0] io_data_12,
  input  [ 7:0] io_data_13,
  input  [ 7:0] io_data_14,
  input  [ 7:0] io_data_15,
  input  [ 7:0] io_data_16,
  input  [ 7:0] io_data_17,
  input  [ 7:0] io_data_18,
  input  [ 7:0] io_data_19,
  input  [ 7:0] io_data_20,
  input  [ 7:0] io_data_21,
  input  [ 7:0] io_data_22,
  input  [ 7:0] io_data_23,
  input  [ 7:0] io_data_24,
  input  [ 7:0] io_data_25,
  input  [ 7:0] io_data_26,
  input  [ 7:0] io_data_27,
  input  [ 7:0] io_data_28,
  input  [ 7:0] io_data_29,
  input  [ 7:0] io_data_30,
  input  [ 7:0] io_data_31,
  input  [ 7:0] io_data_32,
  input  [ 7:0] io_data_33,
  input  [ 7:0] io_data_34,
  input  [ 7:0] io_data_35,
  input  [ 7:0] io_data_36,
  input  [ 7:0] io_data_37,
  input  [ 7:0] io_data_38,
  input  [ 7:0] io_data_39,
  input  [ 7:0] io_data_40,
  input  [ 7:0] io_data_41,
  input  [ 7:0] io_data_42,
  input  [ 7:0] io_data_43,
  input  [ 7:0] io_data_44,
  input  [ 7:0] io_data_45,
  input  [ 7:0] io_data_46,
  input  [ 7:0] io_data_47,
  input  [ 7:0] io_data_48,
  input  [ 7:0] io_data_49,
  input  [ 7:0] io_data_50,
  input  [ 7:0] io_data_51,
  input  [ 7:0] io_data_52,
  input  [ 7:0] io_data_53,
  input  [ 7:0] io_data_54,
  input  [ 7:0] io_data_55,
  input  [ 7:0] io_data_56,
  input  [ 7:0] io_data_57,
  input  [ 7:0] io_data_58,
  input  [ 7:0] io_data_59,
  input  [ 7:0] io_data_60,
  input  [ 7:0] io_data_61,
  input  [ 7:0] io_data_62,
  input  [ 7:0] io_data_63,
  input  [63:0] io_mask,
  input  [ 7:0] io_coreid,
  input  [ 7:0] io_index
);
`ifndef SYNTHESIS
`ifdef DIFFTEST

import "DPI-C" function void v_difftest_SbufferEvent (
  input   longint io_addr,
  input      byte io_data_0,
  input      byte io_data_1,
  input      byte io_data_2,
  input      byte io_data_3,
  input      byte io_data_4,
  input      byte io_data_5,
  input      byte io_data_6,
  input      byte io_data_7,
  input      byte io_data_8,
  input      byte io_data_9,
  input      byte io_data_10,
  input      byte io_data_11,
  input      byte io_data_12,
  input      byte io_data_13,
  input      byte io_data_14,
  input      byte io_data_15,
  input      byte io_data_16,
  input      byte io_data_17,
  input      byte io_data_18,
  input      byte io_data_19,
  input      byte io_data_20,
  input      byte io_data_21,
  input      byte io_data_22,
  input      byte io_data_23,
  input      byte io_data_24,
  input      byte io_data_25,
  input      byte io_data_26,
  input      byte io_data_27,
  input      byte io_data_28,
  input      byte io_data_29,
  input      byte io_data_30,
  input      byte io_data_31,
  input      byte io_data_32,
  input      byte io_data_33,
  input      byte io_data_34,
  input      byte io_data_35,
  input      byte io_data_36,
  input      byte io_data_37,
  input      byte io_data_38,
  input      byte io_data_39,
  input      byte io_data_40,
  input      byte io_data_41,
  input      byte io_data_42,
  input      byte io_data_43,
  input      byte io_data_44,
  input      byte io_data_45,
  input      byte io_data_46,
  input      byte io_data_47,
  input      byte io_data_48,
  input      byte io_data_49,
  input      byte io_data_50,
  input      byte io_data_51,
  input      byte io_data_52,
  input      byte io_data_53,
  input      byte io_data_54,
  input      byte io_data_55,
  input      byte io_data_56,
  input      byte io_data_57,
  input      byte io_data_58,
  input      byte io_data_59,
  input      byte io_data_60,
  input      byte io_data_61,
  input      byte io_data_62,
  input      byte io_data_63,
  input   longint io_mask,
  input      byte io_coreid,
  input      byte io_index
);


  always @(posedge clock) begin
    if (enable)
      v_difftest_SbufferEvent (io_addr, io_data_0, io_data_1, io_data_2, io_data_3, io_data_4, io_data_5, io_data_6, io_data_7, io_data_8, io_data_9, io_data_10, io_data_11, io_data_12, io_data_13, io_data_14, io_data_15, io_data_16, io_data_17, io_data_18, io_data_19, io_data_20, io_data_21, io_data_22, io_data_23, io_data_24, io_data_25, io_data_26, io_data_27, io_data_28, io_data_29, io_data_30, io_data_31, io_data_32, io_data_33, io_data_34, io_data_35, io_data_36, io_data_37, io_data_38, io_data_39, io_data_40, io_data_41, io_data_42, io_data_43, io_data_44, io_data_45, io_data_46, io_data_47, io_data_48, io_data_49, io_data_50, io_data_51, io_data_52, io_data_53, io_data_54, io_data_55, io_data_56, io_data_57, io_data_58, io_data_59, io_data_60, io_data_61, io_data_62, io_data_63, io_mask, io_coreid, io_index);
  end
`endif
`endif
endmodule
