`define LR_RANGE 4:0
`define SRC_RANGE 31:0